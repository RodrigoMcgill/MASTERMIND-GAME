library ieee;
use ieee.std_logic_1164.all;

entity g14_register is
port();

end g14_register;

architecture behavior for g14_register is

begin

end behavior;